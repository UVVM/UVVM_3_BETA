--================================================================================================================================
-- Copyright 2024 UVVM
-- Licensed under the Apache License, Version 2.0 (the "License"); you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at http://www.apache.org/licenses/LICENSE-2.0 and in the provided LICENSE.TXT.
--
-- Unless required by applicable law or agreed to in writing, software distributed under the License is distributed on
-- an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and limitations under the License.
--================================================================================================================================
-- Note : Any functionality not explicitly described in the documentation is subject to change at any time
----------------------------------------------------------------------------------------------------------------------------------

------------------------------------------------------------------------------------------
-- Description   : See library quick reference (under 'doc') and README-file(s)
------------------------------------------------------------------------------------------

context vvc_context is
  library bitvis_vip_axi;
  use bitvis_vip_axi.vvc_transaction_pkg.all;
  use bitvis_vip_axi.vvc_transaction_shared_variables_pkg.all;
  use bitvis_vip_axi.vvc_methods_pkg.all;
  use bitvis_vip_axi.vvc_methods_support_pkg.all;
  use bitvis_vip_axi.vvc_cmd_pkg.all;
  use bitvis_vip_axi.td_vvc_framework_common_methods_pkg.all;
  use bitvis_vip_axi.axi_bfm_pkg.all;
end context;
