--================================================================================================================================
-- Copyright 2020 Bitvis
-- Licensed under the Apache License, Version 2.0 (the "License"); you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at http://www.apache.org/licenses/LICENSE-2.0 and in the provided LICENSE.TXT.
--
-- Unless required by applicable law or agreed to in writing, software distributed under the License is distributed on
-- an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and limitations under the License.
--================================================================================================================================
-- Note : Any functionality not explicitly described in the documentation is subject to change at any time
----------------------------------------------------------------------------------------------------------------------------------

------------------------------------------------------------------------------------------
-- Description   : See library quick reference (under 'doc') and README-file(s)
------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library uvvm_util;
context uvvm_util.uvvm_util_context;

library uvvm_vvc_framework;
use uvvm_vvc_framework.ti_vvc_framework_support_pkg.all;

library bitvis_vip_scoreboard;
use bitvis_vip_scoreboard.generic_sb_support_pkg.all;

library work;
use work.axi_bfm_pkg.all;
use work.axi_channel_handler_pkg.all;
use work.vvc_methods_pkg.all;
use work.vvc_cmd_pkg.all;
use work.td_target_support_pkg.all;
use work.td_vvc_entity_support_pkg.all;
use work.td_cmd_queue_pkg.all;
use work.td_result_queue_pkg.all;
use work.transaction_pkg.all;
use work.axi_read_data_queue_pkg.all;

--=================================================================================================
entity axi_vvc is
    generic(
        GC_ADDR_WIDTH                            : integer range 1 to C_VVC_CMD_ADDR_MAX_LENGTH := 8;
        GC_DATA_WIDTH                            : integer range 1 to C_VVC_CMD_DATA_MAX_LENGTH := 32;
        GC_ID_WIDTH                              : integer range 0 to C_VVC_CMD_ID_MAX_LENGTH   := 8;
        GC_USER_WIDTH                            : integer range 0 to C_VVC_CMD_USER_MAX_LENGTH := 8;
        GC_INSTANCE_IDX                          : natural                                      := 1; -- Instance index for this AXI_VVCT instance
        GC_AXI_CONFIG                            : t_axi_bfm_config                             := C_AXI_BFM_CONFIG_DEFAULT; -- Behavior specification for BFM
        GC_CMD_QUEUE_COUNT_MAX                   : natural                                      := 1000;
        GC_CMD_QUEUE_COUNT_THRESHOLD             : natural                                      := 950;
        GC_CMD_QUEUE_COUNT_THRESHOLD_SEVERITY    : t_alert_level                                := WARNING;
        GC_RESULT_QUEUE_COUNT_MAX                : natural                                      := 1000;
        GC_RESULT_QUEUE_COUNT_THRESHOLD          : natural                                      := 950;
        GC_RESULT_QUEUE_COUNT_THRESHOLD_SEVERITY : t_alert_level                                := WARNING
    );
    port(
        clk               : in    std_logic;
        axi_vvc_master_if : inout t_axi_if := init_axi_if_signals(GC_ADDR_WIDTH, GC_DATA_WIDTH, GC_ID_WIDTH, GC_USER_WIDTH)
    );
begin
    -- Check the interface widths to assure that the interface was correctly set up
    assert (axi_vvc_master_if.write_address_channel.awaddr'length = GC_ADDR_WIDTH) report "axi_vvc_master_if.write_address_channel.awaddr'length =/ GC_ADDR_WIDTH" severity failure;
    assert (axi_vvc_master_if.read_address_channel.araddr'length = GC_ADDR_WIDTH) report "axi_vvc_master_if.read_address_channel.araddr'length =/ GC_ADDR_WIDTH" severity failure;
    assert (axi_vvc_master_if.write_data_channel.wdata'length = GC_DATA_WIDTH) report "axi_vvc_master_if.write_data_channel.wdata'length =/ GC_DATA_WIDTH" severity failure;
    assert (axi_vvc_master_if.write_data_channel.wstrb'length = GC_DATA_WIDTH / 8) report "axi_vvc_master_if.write_data_channel.wstrb'length =/ GC_DATA_WIDTH/8" severity failure;
    assert (axi_vvc_master_if.read_data_channel.rdata'length = GC_DATA_WIDTH) report "axi_vvc_master_if.read_data_channel.rdata'length =/ GC_DATA_WIDTH" severity failure;
end entity axi_vvc;

--=================================================================================================
--=================================================================================================

architecture behave of axi_vvc is

    constant C_SCOPE      : string       := C_VVC_NAME & "," & to_string(GC_INSTANCE_IDX);
    constant C_VVC_LABELS : t_vvc_labels := assign_vvc_labels(C_SCOPE, C_VVC_NAME, GC_INSTANCE_IDX, NA);

    signal executor_is_busy                           : boolean := false;
    signal write_address_channel_executor_is_busy     : boolean := false;
    signal write_data_channel_executor_is_busy        : boolean := false;
    signal write_response_channel_executor_is_busy    : boolean := false;
    signal read_address_channel_executor_is_busy      : boolean := false;
    signal read_data_channel_executor_is_busy         : boolean := false;
    signal any_executors_busy                         : boolean := false;
    signal queue_is_increasing                        : boolean := false;
    signal write_address_channel_queue_is_increasing  : boolean := false;
    signal write_data_channel_queue_is_increasing     : boolean := false;
    signal write_response_channel_queue_is_increasing : boolean := false;
    signal read_address_channel_queue_is_increasing   : boolean := false;
    signal read_data_channel_queue_is_increasing      : boolean := false;
    signal last_cmd_idx_executed                      : natural := natural'high;
    signal last_write_response_channel_idx_executed   : natural := 0;
    signal last_read_data_channel_idx_executed        : natural := 0;
    signal terminate_current_cmd                      : t_flag_record;

    -- Instantiation of the element dedicated Queue
    shared variable command_queue                : work.td_cmd_queue_pkg.t_generic_queue;
    shared variable write_address_channel_queue  : work.td_cmd_queue_pkg.t_generic_queue;
    shared variable write_data_channel_queue     : work.td_cmd_queue_pkg.t_generic_queue;
    shared variable write_response_channel_queue : work.td_cmd_queue_pkg.t_generic_queue;
    shared variable read_address_channel_queue   : work.td_cmd_queue_pkg.t_generic_queue;
    shared variable read_data_channel_queue      : work.td_cmd_queue_pkg.t_generic_queue;
    shared variable result_queue                 : work.td_result_queue_pkg.t_generic_queue;

    -- Transaction info
    alias vvc_transaction_info_trigger        : std_logic is global_axi_vvc_transaction_trigger(GC_INSTANCE_IDX);
    -- VVC Activity
    signal entry_num_in_vvc_activity_register : integer;

    --UVVM: temporary fix for HVVC, remove function below in v3.0
    impure function get_msg_id_panel(   -- v3
        constant command : in t_vvc_cmd_record
    ) return t_msg_id_panel is
    begin
        -- If the parent_msg_id_panel is set then use it,
        -- otherwise use the VVCs msg_id_panel from its config.
        if command.msg(1 to 5) = "HVVC:" then
            return shared_parent_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3
        else
            return shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3
        end if;
    end function;

    impure function queues_are_empty(
        constant void : t_void
    ) return boolean is
        variable v_return : boolean := false;
    begin
        return command_queue.is_empty(VOID) and write_address_channel_queue.is_empty(VOID) and write_data_channel_queue.is_empty(VOID) and write_response_channel_queue.is_empty(VOID) and read_address_channel_queue.is_empty(VOID) and read_data_channel_queue.is_empty(VOID);
    end function;

    impure function get_vvc_config(
        constant void : t_void
    ) return t_vvc_config is
    begin
        return shared_axi_vvc_config.get(GC_INSTANCE_IDX);
    end function get_vvc_config;

    impure function get_vvc_status(
        constant void : t_void
    ) return t_vvc_status is
    begin
        return shared_axi_vvc_status.get(GC_INSTANCE_IDX);
    end function get_vvc_status;

    procedure set_vvc_status(
        constant vvc_status : t_vvc_status
    ) is
    begin
        shared_axi_vvc_status.set(vvc_status, GC_INSTANCE_IDX);
    end procedure set_vvc_status;

    procedure peek_command_and_prepare_executor(
        variable command             : inout t_vvc_cmd_record;
        variable command_queue       : inout work.td_cmd_queue_pkg.t_generic_queue;
        signal   queue_is_increasing : in boolean;
        signal   executor_is_busy    : inout boolean;
        constant vvc_labels          : in t_vvc_labels;
        constant msg_id_panel        : in t_msg_id_panel := shared_msg_id_panel.get(VOID); --UVVM: unused, remove in v3.0
        constant executor_id         : in t_msg_id       := ID_CMD_EXECUTOR;
        constant executor_wait_id    : in t_msg_id       := ID_CMD_EXECUTOR_WAIT
    ) is
        variable v_msg_id_panel : t_msg_id_panel;
        variable v_vvc_status   : t_vvc_status;
    begin
        executor_is_busy              <= false;
        v_vvc_status                  := get_vvc_status(VOID);
        v_vvc_status.previous_cmd_idx := command.cmd_idx;
        v_vvc_status.current_cmd_idx  := 0;
        set_vvc_status(v_vvc_status);

        wait for 0 ns;                  -- to allow delta updates in other processes.
        if command_queue.is_empty(VOID) then
            log(executor_wait_id, "Executor: Waiting for command", to_string(vvc_labels.scope), shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX));
            wait until queue_is_increasing;
        end if;

        -- Queue is now not empty
        executor_is_busy <= true;
        wait until executor_is_busy;
        command          := command_queue.peek(VOID);

        v_msg_id_panel               := get_msg_id_panel(command);
        log(executor_id, to_string(command.proc_call) & " - Will be executed " & format_command_idx(command), to_string(vvc_labels.scope), v_msg_id_panel); -- Get and ack the new command
        v_vvc_status                 := get_vvc_status(VOID);
        v_vvc_status.pending_cmd_cnt := command_queue.get_count(VOID);
        v_vvc_status.current_cmd_idx := command.cmd_idx;
        set_vvc_status(v_vvc_status);
    end procedure peek_command_and_prepare_executor;

begin

    --===============================================================================================
    -- Constructor
    -- - Set up the defaults and show constructor if enabled
    --===============================================================================================
    -- v3
    vvc_constructor(C_SCOPE, GC_INSTANCE_IDX, shared_axi_vvc_config, shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX), command_queue, result_queue, GC_AXI_CONFIG,
                    GC_CMD_QUEUE_COUNT_MAX, GC_CMD_QUEUE_COUNT_THRESHOLD, GC_CMD_QUEUE_COUNT_THRESHOLD_SEVERITY,
                    GC_RESULT_QUEUE_COUNT_MAX, GC_RESULT_QUEUE_COUNT_THRESHOLD, GC_RESULT_QUEUE_COUNT_THRESHOLD_SEVERITY);
    --===============================================================================================

    --===============================================================================================
    -- Set if any of the executors are busy
    --===============================================================================================
    any_executors_busy <= executor_is_busy or write_address_channel_executor_is_busy or write_data_channel_executor_is_busy or write_response_channel_executor_is_busy or read_address_channel_executor_is_busy or read_data_channel_executor_is_busy;
    --===============================================================================================

    --===============================================================================================
    -- Command interpreter
    -- - Interpret, decode and acknowledge commands from the central sequencer
    --===============================================================================================
    cmd_interpreter : process
        variable v_cmd_has_been_acked  : boolean; -- Indicates if acknowledge_cmd() has been called for the current shared_vvc_cmd
        variable v_local_vvc_cmd       : t_vvc_cmd_record := C_VVC_CMD_DEFAULT;
        variable v_msg_id_panel        : t_msg_id_panel;
        variable v_parent_msg_id_panel : t_msg_id_panel; -- v3
        variable v_temp_msg_id_panel   : t_msg_id_panel; --UVVM: temporary fix for HVVC, remove in v3.0
        variable v_vvc_status          : t_vvc_status;
    begin
        -- 0. Initialize the process prior to first command
        work.td_vvc_entity_support_pkg.initialize_interpreter(terminate_current_cmd, global_awaiting_completion);

        -- initialise shared_vvc_last_received_cmd_idx for channel and instance
        shared_vvc_last_received_cmd_idx.set(0, GC_INSTANCE_IDX);

        -- Register VVC in vvc activity register
        entry_num_in_vvc_activity_register <= shared_vvc_activity_register.priv_register_vvc(name                     => C_VVC_NAME,
                                                                                             instance                 => GC_INSTANCE_IDX,
                                                                                             await_selected_supported => false);

        -- Then for every single command from the sequencer
        loop                            -- basically as long as new commands are received

            v_msg_id_panel        := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3
            v_parent_msg_id_panel := get_msg_id_panel(v_local_vvc_cmd); -- v3

            -- 1. wait until command targeted at this VVC. Must match VVC name, instance and channel (if applicable)
            --    releases global semaphore
            -------------------------------------------------------------------------
            work.td_vvc_entity_support_pkg.await_cmd_from_sequencer(C_VVC_LABELS, v_msg_id_panel, v_parent_msg_id_panel, THIS_VVCT, VVC_BROADCAST, global_vvc_busy, global_vvc_ack, v_local_vvc_cmd); -- v3

            v_cmd_has_been_acked := false; -- Clear flag

            -- update shared_vvc_last_received_cmd_idx with received command index
            shared_vvc_last_received_cmd_idx.set(v_local_vvc_cmd.cmd_idx, GC_INSTANCE_IDX);

            -- Select between a provided msg_id_panel via the vvc_cmd_record from a VVC with a higher hierarchy or the
            -- msg_id_panel in this VVC's config. This is to correctly handle the logging when using Hierarchical-VVCs.
            v_msg_id_panel := get_msg_id_panel(v_local_vvc_cmd);

            -- 2a. Put command on the queue if intended for the executor
            -------------------------------------------------------------------------
            if v_local_vvc_cmd.command_type = QUEUED then
                v_vvc_status := get_vvc_status(VOID);
                work.td_vvc_entity_support_pkg.put_command_on_queue(v_local_vvc_cmd, command_queue, v_vvc_status, queue_is_increasing);
                set_vvc_status(v_vvc_status);

            -- 2b. Otherwise command is intended for immediate response
            -------------------------------------------------------------------------
            elsif v_local_vvc_cmd.command_type = IMMEDIATE then

                --UVVM: temporary fix for HVVC, remove two lines below in v3.0
                if v_local_vvc_cmd.operation /= DISABLE_LOG_MSG and v_local_vvc_cmd.operation /= ENABLE_LOG_MSG then
                    v_temp_msg_id_panel := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3
                    shared_axi_vvc_msg_id_panel.set(v_msg_id_panel, GC_INSTANCE_IDX); -- v3         
                end if;

                case v_local_vvc_cmd.operation is

                    when AWAIT_COMPLETION =>
                        work.td_vvc_entity_support_pkg.interpreter_await_completion(v_local_vvc_cmd, command_queue, v_msg_id_panel, any_executors_busy, C_VVC_LABELS, last_cmd_idx_executed); -- v3

                    when AWAIT_ANY_COMPLETION =>
                        if not v_local_vvc_cmd.gen_boolean then
                            -- Called with lastness = NOT_LAST: Acknowledge immediately to let the sequencer continue
                            work.td_target_support_pkg.acknowledge_cmd(global_vvc_ack, v_local_vvc_cmd.cmd_idx);
                            v_cmd_has_been_acked := true;
                        end if;
                        work.td_vvc_entity_support_pkg.interpreter_await_any_completion(v_local_vvc_cmd, command_queue, v_msg_id_panel, any_executors_busy, C_VVC_LABELS, last_cmd_idx_executed, global_awaiting_completion); -- v3

                    when DISABLE_LOG_MSG =>
                        uvvm_util.methods_pkg.disable_log_msg(v_local_vvc_cmd.msg_id, v_msg_id_panel, to_string(v_local_vvc_cmd.msg) & format_command_idx(v_local_vvc_cmd), C_SCOPE, v_local_vvc_cmd.quietness); -- v3

                    when ENABLE_LOG_MSG =>
                        uvvm_util.methods_pkg.enable_log_msg(v_local_vvc_cmd.msg_id, v_msg_id_panel, to_string(v_local_vvc_cmd.msg) & format_command_idx(v_local_vvc_cmd), C_SCOPE, v_local_vvc_cmd.quietness); -- v3

                    when FLUSH_COMMAND_QUEUE =>
                        v_vvc_status := get_vvc_status(VOID);
                        work.td_vvc_entity_support_pkg.interpreter_flush_command_queue(v_local_vvc_cmd, command_queue, v_msg_id_panel, v_vvc_status, C_VVC_LABELS); -- v3
                        work.td_vvc_entity_support_pkg.interpreter_flush_command_queue(v_local_vvc_cmd, write_address_channel_queue, v_msg_id_panel, v_vvc_status, C_VVC_LABELS); -- v3
                        work.td_vvc_entity_support_pkg.interpreter_flush_command_queue(v_local_vvc_cmd, write_data_channel_queue, v_msg_id_panel, v_vvc_status, C_VVC_LABELS); -- v3
                        work.td_vvc_entity_support_pkg.interpreter_flush_command_queue(v_local_vvc_cmd, write_response_channel_queue, v_msg_id_panel, v_vvc_status, C_VVC_LABELS); -- v3
                        work.td_vvc_entity_support_pkg.interpreter_flush_command_queue(v_local_vvc_cmd, read_address_channel_queue, v_msg_id_panel, v_vvc_status, C_VVC_LABELS); -- v3
                        work.td_vvc_entity_support_pkg.interpreter_flush_command_queue(v_local_vvc_cmd, read_data_channel_queue, v_msg_id_panel, v_vvc_status, C_VVC_LABELS); -- v3
                        set_vvc_status(v_vvc_status);

                    when TERMINATE_CURRENT_COMMAND =>
                        work.td_vvc_entity_support_pkg.interpreter_terminate_current_command(v_local_vvc_cmd, v_msg_id_panel, C_VVC_LABELS, terminate_current_cmd); -- v3

                    when FETCH_RESULT =>
                        work.td_vvc_entity_support_pkg.interpreter_fetch_result(result_queue, v_local_vvc_cmd, v_msg_id_panel, C_VVC_LABELS, last_cmd_idx_executed, shared_vvc_response); -- v3

                    when others =>
                        tb_error("Unsupported command received for IMMEDIATE execution: '" & to_string(v_local_vvc_cmd.operation) & "'", C_SCOPE);

                end case;

                --UVVM: temporary fix for HVVC, remove line below in v3.0
                if v_local_vvc_cmd.operation /= DISABLE_LOG_MSG and v_local_vvc_cmd.operation /= ENABLE_LOG_MSG then
                    shared_axi_vvc_msg_id_panel.set(v_temp_msg_id_panel, GC_INSTANCE_IDX); -- v3
                else
                    shared_axi_vvc_msg_id_panel.set(v_msg_id_panel, GC_INSTANCE_IDX); -- v3
                end if;

            else
                tb_error("command_type is not IMMEDIATE or QUEUED", C_SCOPE);
            end if;

            -- 3. Acknowledge command after runing or queuing the command
            -------------------------------------------------------------------------
            if not v_cmd_has_been_acked then
                work.td_target_support_pkg.acknowledge_cmd(global_vvc_ack, v_local_vvc_cmd.cmd_idx);
            end if;

        end loop;
    end process;
    --===============================================================================================

    --===============================================================================================
    -- Updating the activity register
    --===============================================================================================
    p_activity_register_update : process
        variable v_cmd_queues_are_empty : boolean;
    begin
        -- Wait until active and set the activity register to ACTIVE
        if not any_executors_busy then
            wait until any_executors_busy;
        end if;
        v_cmd_queues_are_empty := queues_are_empty(VOID);
        update_vvc_activity_register(global_trigger_vvc_activity_register,
                                     shared_axi_vvc_status,
                                     GC_INSTANCE_IDX,
                                     NA,
                                     ACTIVE,
                                     entry_num_in_vvc_activity_register,
                                     last_cmd_idx_executed,
                                     v_cmd_queues_are_empty,
                                     C_SCOPE);
        -- Wait until inactive and set the activity register to INACTIVE
        if any_executors_busy then
            wait until not any_executors_busy;
        end if;
        v_cmd_queues_are_empty := queues_are_empty(VOID);
        update_vvc_activity_register(global_trigger_vvc_activity_register,
                                     shared_axi_vvc_status,
                                     GC_INSTANCE_IDX,
                                     NA,
                                     INACTIVE,
                                     entry_num_in_vvc_activity_register,
                                     last_cmd_idx_executed,
                                     v_cmd_queues_are_empty,
                                     C_SCOPE);
    end process p_activity_register_update;

    --===============================================================================================
    -- Command executor
    -- - Fetch and execute the commands
    --===============================================================================================
    cmd_executor : process
        variable v_cmd                                   : t_vvc_cmd_record;
        variable v_read_data                             : t_vvc_result; -- See vvc_cmd_pkg
        variable v_timestamp_start_of_current_bfm_access : time                                         := 0 ns;
        variable v_timestamp_start_of_last_bfm_access    : time                                         := 0 ns;
        variable v_timestamp_end_of_last_bfm_access      : time                                         := 0 ns;
        variable v_command_is_bfm_access                 : boolean                                      := false;
        variable v_prev_command_was_bfm_access           : boolean                                      := false;
        variable v_msg_id_panel                          : t_msg_id_panel;
        variable v_normalised_addr                       : unsigned(GC_ADDR_WIDTH - 1 downto 0)         := (others => '0');
        variable v_normalised_data                       : std_logic_vector(GC_DATA_WIDTH - 1 downto 0) := (others => '0');
        variable v_cmd_queues_are_empty                  : boolean;
        variable v_finish2start_warning_triggered        : boolean                                      := false;
        variable v_vvc_config                            : t_vvc_config                                 := get_vvc_config(VOID);
        variable v_vvc_status                            : t_vvc_status;
    begin
        -- 0. Initialize the process prior to first command
        -------------------------------------------------------------------------
        work.td_vvc_entity_support_pkg.initialize_executor(terminate_current_cmd);

        -- Setup AXI scoreboard
        AXI_VVC_SB.set_scope("AXI_VVC_SB");
        AXI_VVC_SB.enable(GC_INSTANCE_IDX, "AXI VVC SB Enabled");
        AXI_VVC_SB.config(GC_INSTANCE_IDX, C_SB_CONFIG_DEFAULT);
        AXI_VVC_SB.enable_log_msg(GC_INSTANCE_IDX, ID_DATA);

        loop

            v_msg_id_panel := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3

            -- 1. Set defaults, fetch command and log
            -------------------------------------------------------------------------
            work.td_vvc_entity_support_pkg.fetch_command_and_prepare_executor(v_cmd, command_queue, v_msg_id_panel, shared_axi_vvc_status, queue_is_increasing, executor_is_busy, C_VVC_LABELS); -- v3

            v_vvc_config := get_vvc_config(VOID);

            -- Select between a provided msg_id_panel via the vvc_cmd_record from a VVC with a higher hierarchy or the
            -- msg_id_panel in this VVC's config. This is to correctly handle the logging when using Hierarchical-VVCs.
            v_msg_id_panel := get_msg_id_panel(v_cmd);

            -- Check if command is a BFM access
            v_prev_command_was_bfm_access := v_command_is_bfm_access; -- save for inter_bfm_delay
            if v_cmd.operation = WRITE or v_cmd.operation = READ or v_cmd.operation = CHECK then
                v_command_is_bfm_access := true;
            else
                v_command_is_bfm_access := false;
            end if;

            -- Insert delay if needed
            work.td_vvc_entity_support_pkg.insert_inter_bfm_delay_if_requested(vvc_config                         => v_vvc_config,
                                                                               command_is_bfm_access              => v_prev_command_was_bfm_access,
                                                                               timestamp_start_of_last_bfm_access => v_timestamp_start_of_last_bfm_access,
                                                                               timestamp_end_of_last_bfm_access   => v_timestamp_end_of_last_bfm_access,
                                                                               msg_id_panel                       => v_msg_id_panel,
                                                                               scope                              => C_SCOPE);

            if v_command_is_bfm_access then
                v_timestamp_start_of_current_bfm_access := now;
            end if;

            -- 2. Execute the fetched command
            -------------------------------------------------------------------------
            case v_cmd.operation is     -- Only operations in the dedicated record are relevant

                -- VVC dedicated operations
                --===================================
                when WRITE =>
                    -- Set vvc transaction info
                    set_global_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);

                    -- Normalise address and data
                    v_normalised_addr := normalize_and_check(v_cmd.addr, v_normalised_addr, ALLOW_WIDER_NARROWER, "v_cmd.addr", "v_normalised_addr", "axi_write() called with to wide address. " & v_cmd.msg);
                    v_normalised_data := normalize_and_check(v_cmd.data_array(0), v_normalised_data, ALLOW_WIDER_NARROWER, "v_cmd.data_array(0)", "v_normalised_data", "axi_write() called with to wide data. " & v_cmd.msg);

                    -- Adding the write command to the write address channel queue , write data channel queue and write response channel queue
                    v_vvc_status := get_vvc_status(VOID);
                    work.td_vvc_entity_support_pkg.put_command_on_queue(v_cmd, write_address_channel_queue, v_vvc_status, write_address_channel_queue_is_increasing);
                    work.td_vvc_entity_support_pkg.put_command_on_queue(v_cmd, write_data_channel_queue, v_vvc_status, write_data_channel_queue_is_increasing);
                    work.td_vvc_entity_support_pkg.put_command_on_queue(v_cmd, write_response_channel_queue, v_vvc_status, write_response_channel_queue_is_increasing);
                    set_vvc_status(v_vvc_status);

                when READ =>
                    -- Set vvc transaction info
                    set_global_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);

                    -- Normalise address and data
                    v_normalised_addr := normalize_and_check(v_cmd.addr, v_normalised_addr, ALLOW_WIDER_NARROWER, "v_cmd.addr", "v_normalised_addr", "axi_read() called with to wide address. " & v_cmd.msg);

                    -- Adding the read command to the read address channel queue and the read address data queue
                    v_vvc_status := get_vvc_status(VOID);
                    work.td_vvc_entity_support_pkg.put_command_on_queue(v_cmd, read_address_channel_queue, v_vvc_status, read_address_channel_queue_is_increasing);
                    work.td_vvc_entity_support_pkg.put_command_on_queue(v_cmd, read_data_channel_queue, v_vvc_status, read_data_channel_queue_is_increasing);
                    set_vvc_status(v_vvc_status);

                when CHECK =>
                    -- Set vvc transaction info
                    set_global_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);

                    -- Normalise address and data
                    v_normalised_addr := normalize_and_check(v_cmd.addr, v_normalised_addr, ALLOW_WIDER_NARROWER, "v_cmd.addr", "v_normalised_addr", "axi_check() called with to wide address. " & v_cmd.msg);
                    v_normalised_data := normalize_and_check(v_cmd.data_array(0), v_normalised_data, ALLOW_WIDER_NARROWER, "v_cmd.data_array(0)", "v_normalised_data", "axi_check() called with to wide data. " & v_cmd.msg);

                    -- Adding the check command to the read address channel queue and the read address data queue
                    v_vvc_status := get_vvc_status(VOID);
                    work.td_vvc_entity_support_pkg.put_command_on_queue(v_cmd, read_address_channel_queue, v_vvc_status, read_address_channel_queue_is_increasing);
                    work.td_vvc_entity_support_pkg.put_command_on_queue(v_cmd, read_data_channel_queue, v_vvc_status, read_data_channel_queue_is_increasing);
                    set_vvc_status(v_vvc_status);

                -- UVVM common operations
                --===================================
                when INSERT_DELAY =>
                    log(ID_INSERTED_DELAY, "Running: " & to_string(v_cmd.proc_call) & " " & format_command_idx(v_cmd), C_SCOPE, v_msg_id_panel);
                    if v_cmd.gen_integer_array(0) = -1 then
                        -- Delay specified using time
                        wait until terminate_current_cmd.is_active = '1' for v_cmd.delay;
                    else
                        -- Delay specified using integer
                        check_value(v_vvc_config.bfm_config.clock_period > -1 ns, TB_ERROR, "Check that clock_period is configured when using insert_delay().",
                                    C_SCOPE, ID_NEVER, v_msg_id_panel);
                        wait until terminate_current_cmd.is_active = '1' for v_cmd.gen_integer_array(0) * v_vvc_config.bfm_config.clock_period;
                    end if;

                when others =>
                    tb_error("Unsupported local command received for execution: '" & to_string(v_cmd.operation) & "'", C_SCOPE);
            end case;

            if v_command_is_bfm_access then
                v_timestamp_end_of_last_bfm_access   := now;
                v_timestamp_start_of_last_bfm_access := v_timestamp_start_of_current_bfm_access;
                if ((v_vvc_config.inter_bfm_delay.delay_type = TIME_START2START) and ((now - v_timestamp_start_of_current_bfm_access) > v_vvc_config.inter_bfm_delay.delay_in_time)) then
                    alert(v_vvc_config.inter_bfm_delay.inter_bfm_delay_violation_severity, "BFM access exceeded specified start-to-start inter-bfm delay, " & to_string(v_vvc_config.inter_bfm_delay.delay_in_time) & ".", C_SCOPE);
                elsif v_vvc_config.inter_bfm_delay.delay_type = TIME_FINISH2START and not v_finish2start_warning_triggered then
                    v_finish2start_warning_triggered := true;
                    tb_warning("Delay type TIME_FINISH2START is not supported by this VVC. Waiting according to TIME_START2START", C_SCOPE);
                end if;
            end if;

            -- Reset terminate flag if any occurred
            if (terminate_current_cmd.is_active = '1') then
                log(ID_CMD_EXECUTOR, "Termination request received", C_SCOPE, v_msg_id_panel);
                uvvm_vvc_framework.ti_vvc_framework_support_pkg.reset_flag(terminate_current_cmd);
            end if;

            -- In case we only allow a single pending transaction, wait here until every channel is finished. 
            -- Even though this wait doesn't have a timeout, each of the executors have timeouts.
            if v_vvc_config.force_single_pending_transaction and v_command_is_bfm_access then
                wait until not write_address_channel_executor_is_busy and not write_data_channel_executor_is_busy and not write_response_channel_executor_is_busy and not read_address_channel_executor_is_busy and not read_data_channel_executor_is_busy;
            end if;

        end loop;
    end process cmd_executor;
    --===============================================================================================

    --===============================================================================================
    -- Read address channel executor
    -- - Fetch and execute the read address channel transactions
    --===============================================================================================
    read_address_channel_executor : process
        variable v_cmd                : t_vvc_cmd_record;
        variable v_msg_id_panel       : t_msg_id_panel;
        variable v_normalized_arid    : std_logic_vector(GC_ID_WIDTH - 1 downto 0) := (others => '0');
        variable v_normalized_araddr  : unsigned(GC_ADDR_WIDTH - 1 downto 0)       := (others => '0');
        variable v_vvc_config         : t_vvc_config                               := get_vvc_config(VOID);
        variable v_vvc_status         : t_vvc_status;
        constant C_CHANNEL_SCOPE      : string                                     := C_VVC_NAME & "_AR" & "," & to_string(GC_INSTANCE_IDX);
        constant C_CHANNEL_VVC_LABELS : t_vvc_labels                               := assign_vvc_labels(C_CHANNEL_SCOPE, C_VVC_NAME, GC_INSTANCE_IDX, NA);

    begin
        -- Set the command response queue up to the same settings as the command queue
        read_address_channel_queue.set_scope(C_CHANNEL_SCOPE & ":Q");
        read_address_channel_queue.set_queue_count_max(v_vvc_config.cmd_queue_count_max);
        read_address_channel_queue.set_queue_count_threshold(v_vvc_config.cmd_queue_count_threshold);
        read_address_channel_queue.set_queue_count_threshold_severity(v_vvc_config.cmd_queue_count_threshold_severity);
        -- Wait until VVC is registered in vvc activity register in the interpreter
        wait until entry_num_in_vvc_activity_register >= 0;

        -- Set initial value of v_msg_id_panel to msg_id_panel in config
        v_msg_id_panel := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3

        loop
            wait for 0 ns;
            -- Fetch commands
            work.td_vvc_entity_support_pkg.fetch_command_and_prepare_executor(v_cmd, read_address_channel_queue, v_msg_id_panel, shared_axi_vvc_status, read_address_channel_queue_is_increasing, read_address_channel_executor_is_busy, C_CHANNEL_VVC_LABELS, ID_CHANNEL_EXECUTOR, ID_CHANNEL_EXECUTOR_WAIT); -- v3

            v_vvc_config := get_vvc_config(VOID);

            -- Select between a provided msg_id_panel via the vvc_cmd_record from a VVC with a higher hierarchy or the
            -- msg_id_panel in this VVC's config. This is to correctly handle the logging when using Hierarchical-VVCs.
            v_msg_id_panel := get_msg_id_panel(v_cmd);

            -- Normalize values from command record to their actual sizes
            if v_normalized_arid'length > 0 then
                v_normalized_arid := normalize_and_check(v_cmd.id, v_normalized_arid, ALLOW_WIDER_NARROWER, "v_cmd.id", "v_normalized_arid", "Function called with to wide arid. " & v_cmd.msg);
            end if;
            v_normalized_araddr := normalize_and_check(v_cmd.addr, v_normalized_araddr, ALLOW_WIDER_NARROWER, "v_cmd.addr", "v_normalized_araddr", "Function called with to araddr. " & v_cmd.msg);
            -- Set vvc transaction info
            set_arw_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);
            -- Start transaction
            read_address_channel_write(arid_value     => v_normalized_arid,
                                       araddr_value   => v_normalized_araddr,
                                       arlen_value    => v_cmd.len,
                                       arsize_value   => v_cmd.size,
                                       arburst_value  => v_cmd.burst,
                                       arlock_value   => v_cmd.lock,
                                       arcache_value  => v_cmd.cache,
                                       arprot_value   => v_cmd.prot,
                                       arqos_value    => v_cmd.qos,
                                       arregion_value => v_cmd.region,
                                       aruser_value   => v_cmd.auser,
                                       msg            => format_msg(v_cmd),
                                       clk            => clk,
                                       arid           => axi_vvc_master_if.read_address_channel.arid,
                                       araddr         => axi_vvc_master_if.read_address_channel.araddr,
                                       arlen          => axi_vvc_master_if.read_address_channel.arlen,
                                       arsize         => axi_vvc_master_if.read_address_channel.arsize,
                                       arburst        => axi_vvc_master_if.read_address_channel.arburst,
                                       arlock         => axi_vvc_master_if.read_address_channel.arlock,
                                       arcache        => axi_vvc_master_if.read_address_channel.arcache,
                                       arprot         => axi_vvc_master_if.read_address_channel.arprot,
                                       arqos          => axi_vvc_master_if.read_address_channel.arqos,
                                       arregion       => axi_vvc_master_if.read_address_channel.arregion,
                                       aruser         => axi_vvc_master_if.read_address_channel.aruser,
                                       arvalid        => axi_vvc_master_if.read_address_channel.arvalid,
                                       arready        => axi_vvc_master_if.read_address_channel.arready,
                                       scope          => C_CHANNEL_SCOPE,
                                       msg_id_panel   => v_msg_id_panel,
                                       config         => v_vvc_config.bfm_config);

            -- Set vvc transaction info back to default values
            reset_arw_vvc_transaction_info(shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd);
        end loop;
    end process read_address_channel_executor;
    --===============================================================================================

    --===============================================================================================
    -- Read data channel executor
    -- - Fetch and execute the read data channel transactions
    --===============================================================================================
    read_data_channel_executor : process
        variable v_cmd                  : t_vvc_cmd_record;
        variable v_result               : t_vvc_result := C_EMPTY_VVC_RESULT; -- See vvc_cmd_pkg
        variable v_msg_id_panel         : t_msg_id_panel;
        variable v_cmd_queues_are_empty : boolean;
        variable v_read_data_queue      : t_axi_read_data_queue;
        variable v_queue_count          : natural;
        variable v_cmd_len              : natural;
        variable v_normalized_rid       : std_logic_vector(GC_ID_WIDTH - 1 downto 0);
        variable v_check_ok             : boolean      := true;
        variable v_vvc_config           : t_vvc_config := get_vvc_config(VOID);
        constant C_CHANNEL_SCOPE        : string       := C_VVC_NAME & "_R" & "," & to_string(GC_INSTANCE_IDX);
        constant C_CHANNEL_VVC_LABELS   : t_vvc_labels := assign_vvc_labels(C_CHANNEL_SCOPE, C_VVC_NAME, GC_INSTANCE_IDX, NA);
    begin
        -- Set the command response queue up to the same settings as the command queue
        read_data_channel_queue.set_scope(C_CHANNEL_SCOPE & ":Q");
        read_data_channel_queue.set_queue_count_max(v_vvc_config.cmd_queue_count_max);
        read_data_channel_queue.set_queue_count_threshold(v_vvc_config.cmd_queue_count_threshold);
        read_data_channel_queue.set_queue_count_threshold_severity(v_vvc_config.cmd_queue_count_threshold_severity);
        -- Setup the read data queue
        v_read_data_queue.set_scope(C_CHANNEL_SCOPE & ":PQ");
        -- Wait until VVC is registered in vvc activity register in the interpreter
        wait until entry_num_in_vvc_activity_register >= 0;

        -- Set initial value of v_msg_id_panel to msg_id_panel in config
        v_msg_id_panel := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3

        loop
            -- get a command from the queue without removing it
            peek_command_and_prepare_executor(v_cmd, read_data_channel_queue, read_data_channel_queue_is_increasing, read_data_channel_executor_is_busy, C_CHANNEL_VVC_LABELS, shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX), ID_CHANNEL_EXECUTOR, ID_CHANNEL_EXECUTOR_WAIT);

            v_vvc_config := get_vvc_config(VOID);

            -- Select between a provided msg_id_panel via the vvc_cmd_record from a VVC with a higher hierarchy or the
            -- msg_id_panel in this VVC's config. This is to correctly handle the logging when using Hierarchical-VVCs.
            v_msg_id_panel := get_msg_id_panel(v_cmd);

            -- Handling commands
            case v_cmd.operation is
                when READ =>
                    -- Set vvc transaction info
                    set_r_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);
                    -- Start transaction
                    read_data_channel_receive(read_result     => v_result,
                                              read_data_queue => v_read_data_queue,
                                              msg             => format_msg(v_cmd),
                                              clk             => clk,
                                              rid             => axi_vvc_master_if.read_data_channel.rid,
                                              rdata           => axi_vvc_master_if.read_data_channel.rdata,
                                              rresp           => axi_vvc_master_if.read_data_channel.rresp,
                                              rlast           => axi_vvc_master_if.read_data_channel.rlast,
                                              ruser           => axi_vvc_master_if.read_data_channel.ruser,
                                              rvalid          => axi_vvc_master_if.read_data_channel.rvalid,
                                              rready          => axi_vvc_master_if.read_data_channel.rready,
                                              scope           => C_CHANNEL_SCOPE,
                                              msg_id_panel    => v_msg_id_panel,
                                              config          => v_vvc_config.bfm_config);

                    -- Looking for the correct response in the queue
                    if v_normalized_rid'length > 0 then
                        v_queue_count := read_data_channel_queue.get_count(VOID);
                        for i in 1 to v_queue_count loop
                            v_cmd            := read_data_channel_queue.peek(POSITION, i);
                            v_normalized_rid := normalize_and_check(v_cmd.id, v_normalized_rid, ALLOW_WIDER_NARROWER, "v_cmd.id", "v_normalized_rid", v_cmd.msg);
                            if check_value(v_result.rid, v_normalized_rid, v_vvc_config.bfm_config.match_strictness, NO_ALERT, "Checking if the correct ID is found in the command queue", C_CHANNEL_SCOPE) then
                                -- Correct ID found. We stop searching for the ID
                                read_data_channel_queue.delete(POSITION, i, SINGLE);
                                exit;
                            elsif i = v_queue_count then
                                -- We didn't find the correct RID
                                error("Unexpected read data with RID: " & to_string(v_result.rid), C_CHANNEL_SCOPE);
                            end if;
                        end loop;
                    else
                        -- ID have length of zero. Using first response in the queue
                        v_cmd := read_data_channel_queue.get(VOID);
                    end if;

                    -- Request SB check result
                    if v_cmd.data_routing = TO_SB then
                        -- call SB check_received
                        AXI_VVC_SB.check_received(GC_INSTANCE_IDX, v_result);
                    else
                        -- Store the result
                        work.td_vvc_entity_support_pkg.store_result(result_queue => result_queue,
                                                                    cmd_idx      => v_cmd.cmd_idx,
                                                                    result       => v_result);
                    end if;

                when CHECK =>
                    -- Set vvc transaction info
                    set_r_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);
                    -- Start transaction
                    read_data_channel_receive(read_result     => v_result,
                                              read_data_queue => v_read_data_queue,
                                              msg             => format_msg(v_cmd),
                                              clk             => clk,
                                              rid             => axi_vvc_master_if.read_data_channel.rid,
                                              rdata           => axi_vvc_master_if.read_data_channel.rdata,
                                              rresp           => axi_vvc_master_if.read_data_channel.rresp,
                                              rlast           => axi_vvc_master_if.read_data_channel.rlast,
                                              ruser           => axi_vvc_master_if.read_data_channel.ruser,
                                              rvalid          => axi_vvc_master_if.read_data_channel.rvalid,
                                              rready          => axi_vvc_master_if.read_data_channel.rready,
                                              scope           => C_CHANNEL_SCOPE,
                                              msg_id_panel    => v_msg_id_panel,
                                              config          => v_vvc_config.bfm_config,
                                              ext_proc_call   => "read_data_channel_check");

                    -- Looking for the correct response in the queue
                    if v_normalized_rid'length > 0 then
                        v_queue_count := read_data_channel_queue.get_count(VOID);
                        for i in 1 to v_queue_count loop
                            v_cmd            := read_data_channel_queue.peek(POSITION, i);
                            v_normalized_rid := normalize_and_check(v_cmd.id, v_normalized_rid, ALLOW_WIDER_NARROWER, "v_cmd.id", "v_normalized_rid", v_cmd.msg);
                            if check_value(v_result.rid, v_normalized_rid, v_vvc_config.bfm_config.match_strictness, NO_ALERT, "Checking if the correct ID is found in the command queue", C_CHANNEL_SCOPE) then
                                -- Correct ID found. We stop searching for the ID
                                read_data_channel_queue.delete(POSITION, i, SINGLE);
                                exit;
                            elsif i = v_queue_count then
                                -- We didn't find the correct RID
                                error("Unexpected read data with RID: " & to_string(v_result.rid), C_CHANNEL_SCOPE);
                            end if;
                        end loop;
                    else
                        -- ID have length of zero. Using first response in the queue
                        v_cmd := read_data_channel_queue.get(VOID);
                    end if;

                    -- Checking response
                    v_cmd_len := to_integer(v_cmd.len);
                    if v_normalized_rid'length > 0 then
                        if not check_value(v_result.rid, v_normalized_rid, v_cmd.alert_level, "Checking RID. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, HEX, SKIP_LEADING_0, ID_POS_ACK, v_msg_id_panel) then
                            v_check_ok := false;
                        end if;
                    end if;
                    if not check_value(v_result.rdata(0 to v_cmd_len), v_cmd.data_array(0 to v_cmd_len), v_cmd.alert_level, "Checking RDATA. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, HEX, SKIP_LEADING_0, ID_POS_ACK, v_msg_id_panel) then
                        v_check_ok := false;
                    end if;
                    if not check_value(v_result.rresp(0 to v_cmd_len) = v_cmd.resp_array(0 to v_cmd_len), v_cmd.alert_level, "Checking RRESP. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, ID_POS_ACK, v_msg_id_panel) then
                        v_check_ok := false;
                    end if;
                    if GC_USER_WIDTH > 0 then
                        if not check_value(v_result.ruser(0 to v_cmd_len), v_cmd.user_array(0 to v_cmd_len), v_cmd.alert_level, "Checking RUSER. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, HEX, SKIP_LEADING_0, ID_POS_ACK, v_msg_id_panel) then
                            v_check_ok := false;
                        end if;
                    end if;

                    if v_check_ok then
                        log(v_vvc_config.bfm_config.id_for_bfm, "read data channel check OK. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, v_msg_id_panel);
                    end if;

                when others =>
                    tb_error("Unsupported local command received for execution: '" & to_string(v_cmd.operation) & "'", C_CHANNEL_SCOPE);
            end case;
            v_check_ok                          := true;
            last_read_data_channel_idx_executed <= v_cmd.cmd_idx;
            -- Set vvc transaction info back to default values
            reset_r_vvc_transaction_info(shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA);
            reset_vvc_transaction_info(shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd);
        end loop;
    end process read_data_channel_executor;
    --===============================================================================================

    --===============================================================================================
    -- write address channel executor
    -- - Fetch and execute the write address channel transactions
    --===============================================================================================
    write_address_channel_executor : process
        variable v_cmd                : t_vvc_cmd_record;
        variable v_msg_id_panel       : t_msg_id_panel;
        variable v_normalized_awid    : std_logic_vector(GC_ID_WIDTH - 1 downto 0) := (others => '0');
        variable v_normalized_awaddr  : unsigned(GC_ADDR_WIDTH - 1 downto 0)       := (others => '0');
        variable v_vvc_config         : t_vvc_config                               := get_vvc_config(VOID);
        constant C_CHANNEL_SCOPE      : string                                     := C_VVC_NAME & "_AW" & "," & to_string(GC_INSTANCE_IDX);
        constant C_CHANNEL_VVC_LABELS : t_vvc_labels                               := assign_vvc_labels(C_CHANNEL_SCOPE, C_VVC_NAME, GC_INSTANCE_IDX, NA);
    begin
        -- Set the command response queue up to the same settings as the command queue
        write_address_channel_queue.set_scope(C_CHANNEL_SCOPE & ":Q");
        write_address_channel_queue.set_queue_count_max(v_vvc_config.cmd_queue_count_max);
        write_address_channel_queue.set_queue_count_threshold(v_vvc_config.cmd_queue_count_threshold);
        write_address_channel_queue.set_queue_count_threshold_severity(v_vvc_config.cmd_queue_count_threshold_severity);

        -- Wait until VVC is registered in vvc activity register in the interpreter
        wait until entry_num_in_vvc_activity_register >= 0;

        -- Set initial value of v_msg_id_panel to msg_id_panel in config
        v_msg_id_panel := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3

        loop
            wait for 0 ns;
            -- Fetch commands
            work.td_vvc_entity_support_pkg.fetch_command_and_prepare_executor(v_cmd, write_address_channel_queue, v_msg_id_panel, shared_axi_vvc_status, write_address_channel_queue_is_increasing, write_address_channel_executor_is_busy, C_CHANNEL_VVC_LABELS, ID_CHANNEL_EXECUTOR, ID_CHANNEL_EXECUTOR_WAIT); -- v3

            v_vvc_config := get_vvc_config(VOID);

            -- Select between a provided msg_id_panel via the vvc_cmd_record from a VVC with a higher hierarchy or the
            -- msg_id_panel in this VVC's config. This is to correctly handle the logging when using Hierarchical-VVCs.
            v_msg_id_panel := get_msg_id_panel(v_cmd);

            -- Normalise address
            if v_normalized_awid'length > 0 then
                v_normalized_awid := normalize_and_check(v_cmd.id, v_normalized_awid, ALLOW_WIDER_NARROWER, "v_cmd.id", "v_normalized_awid", "Function called with to wide awid. " & v_cmd.msg);
            end if;

            v_normalized_awaddr := normalize_and_check(v_cmd.addr, v_normalized_awaddr, ALLOW_WIDER_NARROWER, "v_cmd.addr", "v_normalized_awaddr", "Function called with to awaddr. " & v_cmd.msg);
            -- Set vvc transaction info
            set_arw_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);

            -- Start transaction
            write_address_channel_write(awid_value     => v_normalized_awid,
                                        awaddr_value   => v_normalized_awaddr,
                                        awlen_value    => v_cmd.len,
                                        awsize_value   => v_cmd.size,
                                        awburst_value  => v_cmd.burst,
                                        awlock_value   => v_cmd.lock,
                                        awcache_value  => v_cmd.cache,
                                        awprot_value   => v_cmd.prot,
                                        awqos_value    => v_cmd.qos,
                                        awregion_value => v_cmd.region,
                                        awuser_value   => v_cmd.auser,
                                        msg            => format_msg(v_cmd),
                                        clk            => clk,
                                        awid           => axi_vvc_master_if.write_address_channel.awid,
                                        awaddr         => axi_vvc_master_if.write_address_channel.awaddr,
                                        awlen          => axi_vvc_master_if.write_address_channel.awlen,
                                        awsize         => axi_vvc_master_if.write_address_channel.awsize,
                                        awburst        => axi_vvc_master_if.write_address_channel.awburst,
                                        awlock         => axi_vvc_master_if.write_address_channel.awlock,
                                        awcache        => axi_vvc_master_if.write_address_channel.awcache,
                                        awprot         => axi_vvc_master_if.write_address_channel.awprot,
                                        awqos          => axi_vvc_master_if.write_address_channel.awqos,
                                        awregion       => axi_vvc_master_if.write_address_channel.awregion,
                                        awuser         => axi_vvc_master_if.write_address_channel.awuser,
                                        awvalid        => axi_vvc_master_if.write_address_channel.awvalid,
                                        awready        => axi_vvc_master_if.write_address_channel.awready,
                                        scope          => C_CHANNEL_SCOPE,
                                        msg_id_panel   => v_msg_id_panel,
                                        config         => v_vvc_config.bfm_config);

            -- Set vvc transaction info back to default values
            reset_arw_vvc_transaction_info(shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd);
        end loop;
    end process write_address_channel_executor;
    --===============================================================================================

    --===============================================================================================
    -- write data channel executor
    -- - Fetch and execute the write data channel transactions
    --===============================================================================================
    write_data_channel_executor : process
        variable v_cmd                : t_vvc_cmd_record;
        variable v_msg_id_panel       : t_msg_id_panel;
        variable v_wdata_array_ptr    : t_slv_array_ptr;
        variable v_wstrb_array_ptr    : t_slv_array_ptr;
        variable v_wuser_array_ptr    : t_slv_array_ptr;
        variable v_vvc_config         : t_vvc_config := get_vvc_config(VOID);
        constant C_CHANNEL_SCOPE      : string       := C_VVC_NAME & "_W" & "," & to_string(GC_INSTANCE_IDX);
        constant C_CHANNEL_VVC_LABELS : t_vvc_labels := assign_vvc_labels(C_CHANNEL_SCOPE, C_VVC_NAME, GC_INSTANCE_IDX, NA);
    begin
        -- Set the command response queue up to the same settings as the command queue
        write_data_channel_queue.set_scope(C_CHANNEL_SCOPE & ":Q");
        write_data_channel_queue.set_queue_count_max(v_vvc_config.cmd_queue_count_max);
        write_data_channel_queue.set_queue_count_threshold(v_vvc_config.cmd_queue_count_threshold);
        write_data_channel_queue.set_queue_count_threshold_severity(v_vvc_config.cmd_queue_count_threshold_severity);

        -- Wait until VVC is registered in vvc activity register in the interpreter
        wait until entry_num_in_vvc_activity_register >= 0;

        -- Set initial value of v_msg_id_panel to msg_id_panel in config
        v_msg_id_panel := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3

        loop
            wait for 0 ns;

            -- Fetch commands
            work.td_vvc_entity_support_pkg.fetch_command_and_prepare_executor(v_cmd, write_data_channel_queue, v_msg_id_panel, shared_axi_vvc_status, write_data_channel_queue_is_increasing, write_data_channel_executor_is_busy, C_CHANNEL_VVC_LABELS, ID_CHANNEL_EXECUTOR, ID_CHANNEL_EXECUTOR_WAIT); -- v3

            v_vvc_config := get_vvc_config(VOID);

            -- Select between a provided msg_id_panel via the vvc_cmd_record from a VVC with a higher hierarchy or the
            -- msg_id_panel in this VVC's config. This is to correctly handle the logging when using Hierarchical-VVCs.
            v_msg_id_panel := get_msg_id_panel(v_cmd);

            -- Initializing array pointers
            v_wdata_array_ptr := new t_slv_array(0 to to_integer(unsigned(v_cmd.len)))(GC_DATA_WIDTH-1 downto 0);
            v_wstrb_array_ptr := new t_slv_array(0 to to_integer(unsigned(v_cmd.len)))(GC_DATA_WIDTH/8-1 downto 0);
            v_wuser_array_ptr := new t_slv_array(0 to to_integer(unsigned(v_cmd.len)))(GC_USER_WIDTH-1 downto 0);
            for i in 0 to to_integer(unsigned(v_cmd.len)) loop
                v_wdata_array_ptr(i) := v_cmd.data_array(i)(GC_DATA_WIDTH - 1 downto 0);
                v_wstrb_array_ptr(i) := v_cmd.strb_array(i)(GC_DATA_WIDTH / 8 - 1 downto 0);
                v_wuser_array_ptr(i) := v_cmd.user_array(i)(GC_USER_WIDTH - 1 downto 0);
            end loop;

            -- Set vvc transaction info
            set_w_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);

            -- Start transaction
            write_data_channel_write(wdata_value  => v_wdata_array_ptr.all,
                                     wstrb_value  => v_wstrb_array_ptr.all,
                                     wuser_value  => v_wuser_array_ptr.all,
                                     awlen_value  => v_cmd.len,
                                     msg          => format_msg(v_cmd),
                                     clk          => clk,
                                     wdata        => axi_vvc_master_if.write_data_channel.wdata,
                                     wstrb        => axi_vvc_master_if.write_data_channel.wstrb,
                                     wlast        => axi_vvc_master_if.write_data_channel.wlast,
                                     wuser        => axi_vvc_master_if.write_data_channel.wuser,
                                     wvalid       => axi_vvc_master_if.write_data_channel.wvalid,
                                     wready       => axi_vvc_master_if.write_data_channel.wready,
                                     scope        => C_CHANNEL_SCOPE,
                                     msg_id_panel => v_msg_id_panel,
                                     config       => v_vvc_config.bfm_config);

            deallocate(v_wdata_array_ptr);
            deallocate(v_wstrb_array_ptr);
            deallocate(v_wuser_array_ptr);
            -- Set vvc transaction info back to default values
            reset_w_vvc_transaction_info(shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA);
        end loop;
    end process write_data_channel_executor;
    --===============================================================================================

    --===============================================================================================
    -- write response channel executor
    -- - Fetch and execute the write response channel transactions
    --===============================================================================================
    write_response_channel_executor : process
        variable v_cmd                  : t_vvc_cmd_record;
        variable v_msg_id_panel         : t_msg_id_panel;
        variable v_normalized_bid       : std_logic_vector(GC_ID_WIDTH - 1 downto 0);
        variable v_normalized_buser     : std_logic_vector(GC_USER_WIDTH - 1 downto 0);
        variable v_bid_value            : std_logic_vector(GC_ID_WIDTH - 1 downto 0);
        variable v_bresp_value          : t_xresp;
        variable v_buser_value          : std_logic_vector(GC_USER_WIDTH - 1 downto 0);
        variable v_cmd_queues_are_empty : boolean;
        variable v_queue_count          : integer;
        variable v_vvc_config           : t_vvc_config := get_vvc_config(VOID);
        constant C_CHANNEL_SCOPE        : string       := C_VVC_NAME & "_B" & "," & to_string(GC_INSTANCE_IDX);
        constant C_CHANNEL_VVC_LABELS   : t_vvc_labels := assign_vvc_labels(C_CHANNEL_SCOPE, C_VVC_NAME, GC_INSTANCE_IDX, NA);
    begin
        -- Set the command response queue up to the same settings as the command queue
        write_response_channel_queue.set_scope(C_CHANNEL_SCOPE & ":Q");
        write_response_channel_queue.set_queue_count_max(v_vvc_config.cmd_queue_count_max);
        write_response_channel_queue.set_queue_count_threshold(v_vvc_config.cmd_queue_count_threshold);
        write_response_channel_queue.set_queue_count_threshold_severity(v_vvc_config.cmd_queue_count_threshold_severity);

        -- Wait until VVC is registered in vvc activity register in the interpreter
        wait until entry_num_in_vvc_activity_register >= 0;

        -- Set initial value of v_msg_id_panel to msg_id_panel in config
        v_msg_id_panel := shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX); -- v3

        loop
            -- get a command from the queue without removing it
            peek_command_and_prepare_executor(v_cmd, write_response_channel_queue, write_response_channel_queue_is_increasing, write_response_channel_executor_is_busy, C_CHANNEL_VVC_LABELS, shared_axi_vvc_msg_id_panel.get(GC_INSTANCE_IDX), ID_CHANNEL_EXECUTOR, ID_CHANNEL_EXECUTOR_WAIT);

            v_vvc_config := get_vvc_config(VOID);

            -- Select between a provided msg_id_panel via the vvc_cmd_record from a VVC with a higher hierarchy or the
            -- msg_id_panel in this VVC's config. This is to correctly handle the logging when using Hierarchical-VVCs.
            v_msg_id_panel := get_msg_id_panel(v_cmd);

            -- Set vvc transaction info
            set_b_vvc_transaction_info(vvc_transaction_info_trigger, shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd, v_vvc_config);

            -- Receiving a write response
            write_response_channel_receive(bid_value    => v_bid_value,
                                           bresp_value  => v_bresp_value,
                                           buser_value  => v_buser_value,
                                           msg          => format_msg(v_cmd),
                                           clk          => clk,
                                           bid          => axi_vvc_master_if.write_response_channel.bid,
                                           bresp        => axi_vvc_master_if.write_response_channel.bresp,
                                           buser        => axi_vvc_master_if.write_response_channel.buser,
                                           bvalid       => axi_vvc_master_if.write_response_channel.bvalid,
                                           bready       => axi_vvc_master_if.write_response_channel.bready,
                                           alert_level  => error,
                                           scope        => C_CHANNEL_SCOPE,
                                           msg_id_panel => v_msg_id_panel,
                                           config       => v_vvc_config.bfm_config);

            -- Looking for the correct response in the queue
            if v_normalized_bid'length > 0 then
                v_queue_count := write_response_channel_queue.get_count(VOID);
                for i in 1 to v_queue_count loop
                    v_cmd            := write_response_channel_queue.peek(POSITION, i);
                    v_normalized_bid := normalize_and_check(v_cmd.id, v_normalized_bid, ALLOW_WIDER_NARROWER, "v_cmd.id", "v_normalized_bid", v_cmd.msg);
                    if check_value(v_bid_value, v_normalized_bid, v_vvc_config.bfm_config.match_strictness, NO_ALERT, "Checking if the correct ID is found in the command queue", C_CHANNEL_SCOPE) then
                        -- Correct ID found. We stop searching for the ID
                        write_response_channel_queue.delete(POSITION, i, SINGLE);
                        exit;
                    elsif i = v_queue_count then
                        -- We didn't find the correct BID
                        error("Unexpected write response with BID: " & to_string(v_bid_value), C_CHANNEL_SCOPE);
                    end if;
                end loop;
            else
                -- ID have length of zero. Using first response in the queue
                v_cmd := write_response_channel_queue.get(VOID);
            end if;

            -- Checking response
            if v_normalized_bid'length > 0 then
                check_value(v_bid_value, v_normalized_bid, v_vvc_config.bfm_config.match_strictness, error, "Checking BID value. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, HEX, KEEP_LEADING_0, ID_POS_ACK, v_msg_id_panel);
            end if;
            if v_normalized_buser'length > 0 then
                v_normalized_buser := normalize_and_check(v_cmd.user, v_normalized_buser, ALLOW_WIDER_NARROWER, "v_cmd.user", "v_normalized_buser", v_cmd.msg);
                check_value(v_buser_value, v_normalized_buser, v_vvc_config.bfm_config.match_strictness, error, "Checking BUSER value. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, HEX, KEEP_LEADING_0, ID_POS_ACK, v_msg_id_panel);
            end if;
            check_value(v_bresp_value = v_cmd.resp, error, "Checking BRESP value. " & add_msg_delimiter(format_msg(v_cmd)), C_CHANNEL_SCOPE, ID_POS_ACK, v_msg_id_panel);

            last_write_response_channel_idx_executed <= v_cmd.cmd_idx;
            -- Set vvc transaction info back to default values
            reset_b_vvc_transaction_info(shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA);
            reset_vvc_transaction_info(shared_axi_vvc_transaction_info, GC_INSTANCE_IDX, NA, v_cmd);
        end loop;
    end process write_response_channel_executor;
    --===============================================================================================

    --===============================================================================================
    -- Command termination handler
    -- - Handles the termination request record (sets and resets terminate flag on request)
    --===============================================================================================
    cmd_terminator : uvvm_vvc_framework.ti_vvc_framework_support_pkg.flag_handler(terminate_current_cmd); -- flag: is_active, set, reset
    --===============================================================================================

end architecture behave;
